
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
ENTITY full_adder_tb IS
END full_adder_tb;
 
ARCHITECTURE full_adder_testbench OF  full_adder_tb IS
 

 
COMPONENT full_adder is
 PORT(
 A : IN std_logic;
 B : IN std_logic;
 Cin : IN std_logic;
 S : OUT std_logic;
 Cout : OUT std_logic
 );
END COMPONENT;
 
signal A : std_logic := '0';
signal B : std_logic := '0';
signal Cin : std_logic := '0';
 
signal S : std_logic;
signal Cout : std_logic;
 
BEGIN
 

 uut: full_adder
 PORT MAP (
 A => A,
 B => B,
 Cin => Cin,
 S => S,
 Cout => Cout
 );
 

 process
 begin
 
  wait for 10 ns;
 

  A <= '1';
  B <= '0';
  Cin <= '0';
  wait for 10 ns;
  
  A <= '0';
  B <= '1';
  Cin <= '0';
  wait for 10 ns;
 
  A <= '1';
  B <= '1';
  Cin <= '0';
  wait for 10 ns;
 
  A <= '0';
  B <= '0';
  Cin <= '1';
  wait for 10 ns;
 
  A <= '1';
  B <= '0';
  Cin <= '1';
  wait for 10 ns;
 
  A <= '0';
  B <= '1';
  Cin <= '1';
  wait for 10 ns;
 
  A <= '1';
  B <= '1';
  Cin <= '1';
  wait for 10 ns;
  
  WAIT;
 
 end process;
 
END full_adder_testbench;

